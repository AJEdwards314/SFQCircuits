.subckt DCSFQ 2 17
B01        5          3          jj1     area=1.32
B02        5          6          jj1     area=1
B03        9          10         jj1     area=1.5
B04        13         14         jj1     area=1.96
B05        15         16         jj1     area=1.96
IB01       0          8          pwl(0 0 5p 162.5u)
IB02       0          12         pwl(0 0 5p 260u)
L01        2          1          0.848p
L02        0          1          7.712p
L03        1          3          1.778p
L04        5          7          0.543p
L05        7          9          3.149p
L06        9          11         1.323p
L07        11         13         1.095p
L08        13         15         2.951p
L09        15         17         1.63p
LP01       0          6          0.398p
LP02       0          10         0.211p
LP03       0          14         0.276p
LP04       0          16         0.224p
LPR01      7          8          0.915p
LPR02      11         12         0.307p
LRB01      4          5          1p
LRB02      18         6          1p
LRB03      19         10         1p
LRB04      20         14         1p
LRB05      21         16         1p
RB01       3          4          8.56
RB02       18         5          11.30
RB03       19         9          7.53
RB04       20         13         5.77
RB05       21         15         5.77
.model jj1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.ends DCSFQ

.subckt CONFLU 1 2 3 4 14
B01 5 0 jmitll
B02 5 9 jmitll area=1.5
B03 6 0 jmitll
B04 6 10 jmitll area=1.5
B05 7 0 jmitll
B06 7 11 jmitll area=1.5
B07 8 0 jmitll
B08 8 12 jmitll area=1.5
B0L 14 0 jmitll
L01 1 5 0.5p
L02 2 6 0.5p
L03 3 7 0.5p
L04 4 8 0.5p
L05 9 13 0.5p
L06 10 13 0.5p
L07 11 13 0.5p
L08 12 13 0.5p
LC1 13 14 2p
I01 0 13 pwl(0 0 5p 800u)
.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.ends CONFLU

.subckt NEURON 11 5 4
B01        0          11         jmitll
B02        0          4          jmitll
B03        0          5          jmitll
IB0        0          11         pwl(0 0 5p 0u)
L02        11         2          5p
L03        5          6          5p
L04        3          4          5p
K01        L04        L03        0.6
R01        2          3          0.5
R02        3          0          0.075
R03        6          0          0.2
.ends NEURON

.subckt SYNAPSE 1 9
B01        7          2          jmitll
B02        0          7          jmitll
IB0        0          6          pwl(0 0 5p 100u)
L01        7          9          0.1p
L02        6          7          0.1p
R0L        9          0          1
X01 DCSFQ  1          2
.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.ends SYNAPSE

.subckt SYNEURON 1 2 4
X01 NEURON 1 2 3
X02 SYNAPSE 3 4
.ends SYNEURON

.subckt SPLITTER 1 11 10
# Junctions
B01	2	0	 jmitll
B02	4	0	 jmitll
B03	5	0	 jmitll
B04	6	0	 jmitll
B05	7	0	 jmitll
B06	6	8	 jmitll2
B07	7	9	 jmitll2

# Inductors
L01	1	2	0.5p
L02	2	3	0.5p
L03	3	5	0.5p
L04	3	4	0.5p
L05	5	7	0.5p
L06	4	6	0.5p
L07	9	11	0.5p
L08	8	10	0.5p

# Bias Currents
I01	3	0	 pwl(0 0 5p 250u)
I02	9	0	 pwl(0 0 5p 175u)
I03	8	0	 pwl(0 0 5p 175u)

# Resistors
R0L1    11  0   1
R0L2    10  0   1
R0L     3   0   1
.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.2mA)
.model jmitll2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.1mA)
.ends SPLITTER