* Synaptic Test Circuit 

.SUBCKT DCSFQ 2 17
B01        5          3          jj1 area=1.5
B02        5          6          jj1  
B03        9          10         jj1     
B04        13         14         jj1     
B05        15         16         jj1 
IB01       0          8          pwl(0 0 5p 30u)
IB02       0          12         pwl(0 0 5p 300u)
L03        2          3          1p    
L04        5          7          0.5p    
L05        7          9          3p    
L06        9          11         1p    
L07        11         13         1p    
L08        13         15         3p    
L09        15         17         0.1p     
LP01       0          6          0.1p    
LP02       0          10         0.1p    
LP03       0          14         0.1p    
LP04       0          16         0.1p    
LPR01      7          8          0.1p    
LPR02      11         12         0.1p    
LRB01      4          5          0.5p        
LRB02      18         6          0.5p        
LRB03      19         10         0.5p        
LRB04      20         14         0.5p        
LRB05      21         16         0.5p             
RB03       19         9          6   
RB04       20         13         8
RB05       21         15         6
.model jj1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.1mA)
.ends DCSFQ

B01        7          2          jmitll     
B02        0          7          jmitll     
IB0        0          6          pwl(0 0 5p 100u)
L01        7          9          0.1p    
L02        6          7          0.1p 
R0L        9          0          1
X01 DCSFQ  1          2
Vin	1	0   pulse(0 450u 0 4.5952p 4.5952p 0 20p)

.temp 0
.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.tran 0.005p 100p 0 0.005p 
.print DEVV VIN 
.print PHASE B01 
.print PHASE B02
.print NODEV 2 0
.print NODEV 9 0
.end