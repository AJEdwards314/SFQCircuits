.subckt DCSFQ 2 17
B01        5          3          jj1     area=1.32
B02        5          6          jj1     area=1
B03        9          10         jj1     area=1.5
B04        13         14         jj1     area=1.96
B05        15         16         jj1     area=1.96
IB01       0          8          pwl(0 0 5p 162.5u)
IB02       0          12         pwl(0 0 5p 260u)
L01        2          1          0.848p
L02        0          1          7.712p
L03        1          3          1.778p
L04        5          7          0.543p
L05        7          9          3.149p
L06        9          11         1.323p
L07        11         13         1.095p
L08        13         15         2.951p
L09        15         17         1.63p
LP01       0          6          0.398p
LP02       0          10         0.211p
LP03       0          14         0.276p
LP04       0          16         0.224p
LPR01      7          8          0.915p
LPR02      11         12         0.307p
LRB01      4          5          1p
LRB02      18         6          1p
LRB03      19         10         1p
LRB04      20         14         1p
LRB05      21         16         1p
RB01       3          4          8.56
RB02       18         5          11.30
RB03       19         9          7.53
RB04       20         13         5.77
RB05       21         15         5.77
.model jj1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.ends DCSFQ

.subckt CONFLU 1 2 3 4 14
B01 5 0 jmitll
B02 5 9 jmitll area=1.5
B03 6 0 jmitll
B04 6 10 jmitll area=1.5
B05 7 0 jmitll
B06 7 11 jmitll area=1.5
B07 8 0 jmitll
B08 8 12 jmitll area=1.5
B0L 14 0 jmitll
L01 1 5 0.5p
L02 2 6 0.5p
L03 3 7 0.5p
L04 4 8 0.5p
L05 9 13 0.5p
L06 10 13 0.5p
L07 11 13 0.5p
L08 12 13 0.5p
LC1 13 14 2p
I01 0 13 pwl(0 0 5p 800u)
.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.ends CONFLU

.subckt NEURON 11 5 4
B01        0          11         jmitll
B02        0          4          jmitll
B03        0          5          jmitll
IB0        0          11         pwl(0 0 5p 0u)
L02        11         2          5p
L03        5          6          5p
L04        3          4          5p
K01        L04        L03        0.6
R01        2          3          0.5
R02        3          0          0.075
R03        6          0          0.2
.ends NEURON

.subckt SYNAPSE 1 6 9
B01        7          2          jmitll
B02        0          7          jmitll
L01        7          9          0.1p
L02        6          7          0.1p
R0L        9          0          1
X01 DCSFQ  1          2
.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.ends SYNAPSE

.subckt SPLITTER 1 11 10
# Junctions
B01	2	0	 jmitll
B02	4	0	 jmitll
B03	5	0	 jmitll
B04	6	0	 jmitll
B05	7	0	 jmitll
B06	6	8	 jmitll2
B07	7	9	 jmitll2

# Inductors
L01	1	2	0.5p
L02	2	3	0.5p
L03	3	5	0.5p
L04	3	4	0.5p
L05	5	7	0.5p
L06	4	6	0.5p
L07	9	11	0.5p
L08	8	10	0.5p

# Bias Currents
I01	3	0	 pwl(0 0 5p 250u)
I02	9	0	 pwl(0 0 5p 175u)
I03	8	0	 pwl(0 0 5p 175u)

# Resistors
R0L1    11  0   1
R0L2    10  0   1
R0L     3   0   1
.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.2mA)
.model jmitll2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.1mA)
.ends SPLITTER
VIN1 1 0 pwl(0 0 1.9477548542880714e-11 0 2.4477548542880713e-11 0.00041 2.9477548542880715e-11 0 5.618304419565179e-11 0 6.118304419565179e-11 0.00041 6.618304419565179e-11 0 5.6896084048857785e-11 0 6.189608404885779e-11 0.00041 6.689608404885778e-11 0 5.6977779809382e-11 0 6.1977779809382e-11 0.00041 6.6977779809382e-11 0 7.679012322438772e-11 0 8.179012322438772e-11 0.00041 8.679012322438771e-11 0 1.354679788720895e-10 0 1.404679788720895e-10 0.00041 1.4546797887208951e-10 0 1.5971696516810982e-10 0 1.6471696516810983e-10 0.00041 1.6971696516810984e-10 0 1.8690781404982388e-10 0 1.9190781404982388e-10 0.00041 1.969078140498239e-10 0 2.883121092965499e-10 0 2.9331210929654987e-10 0.00041 2.9831210929654986e-10 0 5.063912201924822e-10 0 5.113912201924822e-10 0.00041 5.163912201924822e-10 0 6.247026374766568e-10 0 6.297026374766568e-10 0.00041 6.347026374766568e-10 0 6.247489964887105e-10 0 6.297489964887104e-10 0.00041 6.347489964887104e-10 0 7.064364044023191e-10 0 7.114364044023191e-10 0.00041 7.164364044023191e-10 0 )
VIN2 2 0 pwl(0 0 6.6559754966098765e-12 0 1.1655975496609876e-11 0.00041 1.6655975496609875e-11 0 2.413478295031041e-11 0 2.913478295031041e-11 0.00041 3.413478295031041e-11 0 2.447432573755136e-11 0 2.947432573755136e-11 0.00041 3.447432573755136e-11 0 2.451322848065813e-11 0 2.951322848065813e-11 0.00041 3.451322848065813e-11 0 3.394767772589895e-11 0 3.894767772589895e-11 0.00041 4.3947677725898955e-11 0 6.188951374861412e-11 0 6.688951374861412e-11 0.00041 7.188951374861411e-11 0 7.343665008005238e-11 0 7.843665008005238e-11 0.00041 8.343665008005237e-11 0 8.638467335705908e-11 0 9.138467335705908e-11 0.00041 9.638467335705907e-11 0 1.346724329983572e-10 0 1.3967243299835722e-10 0.00041 1.4467243299835722e-10 0 2.3851962866308704e-10 0 2.43519628663087e-10 0.00041 2.48519628663087e-10 0 2.9485839879840835e-10 0 2.9985839879840833e-10 0.00041 3.048583987984083e-10 0 2.9488047451843387e-10 0 2.9988047451843385e-10 0.00041 3.0488047451843383e-10 0 3.3377924019158086e-10 0 3.3877924019158084e-10 0.00041 3.437792401915808e-10 0 3.350220576473504e-10 0 3.400220576473504e-10 0.00041 3.4502205764735036e-10 0 3.53354634255933e-10 0 3.5835463425593297e-10 0.00041 3.6335463425593296e-10 0 3.679077719052679e-10 0 3.729077719052679e-10 0.00041 3.779077719052679e-10 0 4.219062059522135e-10 0 4.269062059522135e-10 0.00041 4.3190620595221347e-10 0 4.279749495326692e-10 0 4.329749495326692e-10 0.00041 4.379749495326692e-10 0 4.33239711926298e-10 0 4.3823971192629797e-10 0.00041 4.4323971192629795e-10 0 4.588206161513155e-10 0 4.638206161513155e-10 0.00041 4.688206161513155e-10 0 4.594549738447844e-10 0 4.644549738447844e-10 0.00041 4.694549738447844e-10 0 4.6177493062565087e-10 0 4.667749306256508e-10 0.00041 4.717749306256508e-10 0 4.794354695968356e-10 0 4.844354695968356e-10 0.00041 4.894354695968356e-10 0 4.927134390478047e-10 0 4.977134390478046e-10 0.00041 5.027134390478046e-10 0 5.225022135056444e-10 0 5.275022135056444e-10 0.00041 5.325022135056444e-10 0 5.295937006913822e-10 0 5.345937006913822e-10 0.00041 5.395937006913822e-10 0 5.372773137773502e-10 0 5.422773137773502e-10 0.00041 5.472773137773502e-10 0 5.690274683998695e-10 0 5.740274683998695e-10 0.00041 5.790274683998695e-10 0 5.986025588591212e-10 0 6.036025588591212e-10 0.00041 6.086025588591211e-10 0 6.041475749771314e-10 0 6.091475749771314e-10 0.00041 6.141475749771314e-10 0 6.077606279064736e-10 0 6.127606279064736e-10 0.00041 6.177606279064736e-10 0 6.287313815025132e-10 0 6.337313815025132e-10 0.00041 6.387313815025132e-10 0 6.379597964157198e-10 0 6.429597964157198e-10 0.00041 6.479597964157197e-10 0 6.526115408794459e-10 0 6.576115408794459e-10 0.00041 6.626115408794459e-10 0 )
VIN3 3 0 pwl(0 0 3.961598233416525e-10 0 4.0115982334165247e-10 0.00041 4.0615982334165245e-10 0 9.977221132065063e-10 0 1.0027221132065064e-09 0.00041 1.0077221132065065e-09 0 )
VIN4 4 0 pwl(0 0 3.5795914238134605e-11 0 4.079591423813461e-11 0.00041 4.579591423813461e-11 0 9.697174032608654e-11 0 1.0197174032608653e-10 0.00041 1.0697174032608653e-10 0 9.816014008142986e-11 0 1.0316014008142986e-10 0.00041 1.0816014008142985e-10 0 9.829629968230355e-11 0 1.0329629968230354e-10 0.00041 1.0829629968230354e-10 0 1.3131687204064646e-10 0 1.3631687204064647e-10 0.00041 1.4131687204064648e-10 0 2.291132981201497e-10 0 2.341132981201497e-10 0.00041 2.391132981201497e-10 0 2.6952827528018367e-10 0 2.7452827528018365e-10 0.00041 2.7952827528018363e-10 0 3.148463567497072e-10 0 3.1984635674970716e-10 0.00041 3.2484635674970715e-10 0 4.838535154942508e-10 0 4.888535154942508e-10 0.00041 4.938535154942508e-10 0 8.473187003208055e-10 0 8.523187003208055e-10 0.00041 8.573187003208054e-10 0 )
VIN5 5 0 pwl(0 0 1.7993190396890958e-12 0 6.7993190396890955e-12 0.00041 1.1799319039689095e-11 0 1.1995290054347743e-11 0 1.6995290054347742e-11 0.00041 2.199529005434774e-11 0 1.2193356680238297e-11 0 1.7193356680238296e-11 0.00041 2.2193356680238295e-11 0 1.2216049947050578e-11 0 1.7216049947050577e-11 0.00041 2.2216049947050576e-11 0 1.771947867344106e-11 0 2.271947867344106e-11 0.00041 2.7719478673441058e-11 0 3.401888302002491e-11 0 3.901888302002491e-11 0.00041 4.4018883020024913e-11 0 4.0754712546697226e-11 0 4.575471254669723e-11 0.00041 5.075471254669723e-11 0 4.8307726124951136e-11 0 5.330772612495114e-11 0.00041 5.830772612495113e-11 0 7.64755859157084e-11 0 8.147558591570839e-11 0.00041 8.647558591570839e-11 0 1.370531167201341e-10 0 1.4205311672013412e-10 0.00041 1.4705311672013412e-10 0 1.6991739929907154e-10 0 1.7491739929907155e-10 0.00041 1.7991739929907156e-10 0 1.6993027680241977e-10 0 1.7493027680241978e-10 0.00041 1.7993027680241979e-10 0 1.9262122344508884e-10 0 1.9762122344508885e-10 0.00041 2.0262122344508886e-10 0 1.9334620029428777e-10 0 1.9834620029428777e-10 0.00041 2.0334620029428778e-10 0 2.0404020331596094e-10 0 2.0904020331596095e-10 0.00041 2.1404020331596096e-10 0 2.125295336114063e-10 0 2.1752953361140632e-10 0.00041 2.2252953361140632e-10 0 2.440286201387913e-10 0 2.4902862013879126e-10 0.00041 2.5402862013879124e-10 0 2.4756872056072375e-10 0 2.5256872056072374e-10 0.00041 2.575687205607237e-10 0 2.506398319570072e-10 0 2.556398319570072e-10 0.00041 2.606398319570072e-10 0 2.6556202608826744e-10 0 2.705620260882674e-10 0.00041 2.755620260882674e-10 0 2.659320680761243e-10 0 2.709320680761243e-10 0.00041 2.7593206807612427e-10 0 2.6728537619829637e-10 0 2.7228537619829635e-10 0.00041 2.7728537619829634e-10 0 2.775873572648208e-10 0 2.825873572648208e-10 0.00041 2.8758735726482077e-10 0 2.853328394445528e-10 0 2.9033283944455277e-10 0.00041 2.9533283944455276e-10 0 3.0270962454495933e-10 0 3.077096245449593e-10 0.00041 3.127096245449593e-10 0 3.068463254033064e-10 0 3.1184632540330636e-10 0.00041 3.1684632540330635e-10 0 3.113284330367877e-10 0 3.1632843303678767e-10 0.00041 3.2132843303678765e-10 0 3.298493565665906e-10 0 3.348493565665906e-10 0.00041 3.398493565665906e-10 0 3.4710149266782073e-10 0 3.521014926678207e-10 0.00041 3.571014926678207e-10 0 3.503360854033267e-10 0 3.5533608540332667e-10 0.00041 3.6033608540332665e-10 0 3.524436996121096e-10 0 3.5744369961210957e-10 0.00041 3.6244369961210956e-10 0 3.646766392097994e-10 0 3.6967663920979936e-10 0.00041 3.7467663920979934e-10 0 3.700598812425032e-10 0 3.7505988124250317e-10 0.00041 3.8005988124250315e-10 0 3.786067321796768e-10 0 3.836067321796768e-10 0.00041 3.886067321796768e-10 0 3.8909395428237484e-10 0 3.9409395428237483e-10 0.00041 3.990939542823748e-10 0 4.0141566072135247e-10 0 4.0641566072135245e-10 0.00041 4.1141566072135243e-10 0 4.306973538544831e-10 0 4.356973538544831e-10 0.00041 4.4069735385448306e-10 0 4.322342414403645e-10 0 4.372342414403645e-10 0.00041 4.422342414403645e-10 0 4.468922905922227e-10 0 4.518922905922227e-10 0.00041 4.568922905922227e-10 0 4.581346658829152e-10 0 4.631346658829152e-10 0.00041 4.681346658829152e-10 0 4.771151700662107e-10 0 4.821151700662107e-10 0.00041 4.871151700662107e-10 0 4.831050898076728e-10 0 4.881050898076728e-10 0.00041 4.931050898076728e-10 0 4.877919364508718e-10 0 4.927919364508717e-10 0.00041 4.977919364508717e-10 0 4.959630096156474e-10 0 5.009630096156474e-10 0.00041 5.059630096156474e-10 0 4.986077023991868e-10 0 5.036077023991868e-10 0.00041 5.086077023991868e-10 0 5.06065927289239e-10 0 5.11065927289239e-10 0.00041 5.16065927289239e-10 0 5.071265478490253e-10 0 5.121265478490253e-10 0.00041 5.171265478490253e-10 0 5.235960217857286e-10 0 5.285960217857285e-10 0.00041 5.335960217857285e-10 0 5.463884034615215e-10 0 5.513884034615215e-10 0.00041 5.563884034615215e-10 0 5.519094282069006e-10 0 5.569094282069006e-10 0.00041 5.619094282069005e-10 0 5.835367377340053e-10 0 5.885367377340053e-10 0.00041 5.935367377340053e-10 0 5.846137640484927e-10 0 5.896137640484927e-10 0.00041 5.946137640484927e-10 0 5.874091919557479e-10 0 5.924091919557479e-10 0.00041 5.974091919557479e-10 0 5.903816787860721e-10 0 5.953816787860721e-10 0.00041 6.003816787860721e-10 0 5.980172481553577e-10 0 6.030172481553577e-10 0.00041 6.080172481553576e-10 0 6.07374700760351e-10 0 6.12374700760351e-10 0.00041 6.17374700760351e-10 0 6.127341288681853e-10 0 6.177341288681853e-10 0.00041 6.227341288681853e-10 0 6.139796692092079e-10 0 6.189796692092078e-10 0.00041 6.239796692092078e-10 0 6.339595827749054e-10 0 6.389595827749054e-10 0.00041 6.439595827749054e-10 0 6.389342219294889e-10 0 6.439342219294889e-10 0.00041 6.489342219294889e-10 0 6.400699210760943e-10 0 6.450699210760942e-10 0.00041 6.500699210760942e-10 0 6.477822853514718e-10 0 6.527822853514718e-10 0.00041 6.577822853514718e-10 0 )
X6 SPLITTER 1 6 7
X7 SPLITTER 7 8 9
X8 SPLITTER 2 10 11
X9 SPLITTER 11 12 13
X10 SPLITTER 3 14 15
X11 SPLITTER 15 16 17
X12 SPLITTER 4 18 19
X13 SPLITTER 19 20 21
IB22 6 0 pwl(0 0 5p 118.642u)
X23 SYNAPSE 6 0 23
IB24 10 0 pwl(0 0 5p 120.474u)
X25 SYNAPSE 0 10 25
IB27 14 0 pwl(0 0 5p 118.762u)
X28 SYNAPSE 14 0 28
IB29 18 0 pwl(0 0 5p 127.69u)
X30 SYNAPSE 18 0 30
IB31 31 0 pwl(0 0 5p 116.798u)
VIN31 31 0 pwl(0 0 1.7993190396890958e-12 0 6.7993190396890955e-12 0.00041 1.1799319039689095e-11 0 1.1995290054347743e-11 0 1.6995290054347742e-11 0.00041 2.199529005434774e-11 0 1.2193356680238297e-11 0 1.7193356680238296e-11 0.00041 2.2193356680238295e-11 0 1.2216049947050578e-11 0 1.7216049947050577e-11 0.00041 2.2216049947050576e-11 0 1.771947867344106e-11 0 2.271947867344106e-11 0.00041 2.7719478673441058e-11 0 3.401888302002491e-11 0 3.901888302002491e-11 0.00041 4.4018883020024913e-11 0 4.0754712546697226e-11 0 4.575471254669723e-11 0.00041 5.075471254669723e-11 0 4.8307726124951136e-11 0 5.330772612495114e-11 0.00041 5.830772612495113e-11 0 7.64755859157084e-11 0 8.147558591570839e-11 0.00041 8.647558591570839e-11 0 1.370531167201341e-10 0 1.4205311672013412e-10 0.00041 1.4705311672013412e-10 0 1.6991739929907154e-10 0 1.7491739929907155e-10 0.00041 1.7991739929907156e-10 0 1.6993027680241977e-10 0 1.7493027680241978e-10 0.00041 1.7993027680241979e-10 0 1.9262122344508884e-10 0 1.9762122344508885e-10 0.00041 2.0262122344508886e-10 0 1.9334620029428777e-10 0 1.9834620029428777e-10 0.00041 2.0334620029428778e-10 0 2.0404020331596094e-10 0 2.0904020331596095e-10 0.00041 2.1404020331596096e-10 0 2.125295336114063e-10 0 2.1752953361140632e-10 0.00041 2.2252953361140632e-10 0 2.440286201387913e-10 0 2.4902862013879126e-10 0.00041 2.5402862013879124e-10 0 2.4756872056072375e-10 0 2.5256872056072374e-10 0.00041 2.575687205607237e-10 0 2.506398319570072e-10 0 2.556398319570072e-10 0.00041 2.606398319570072e-10 0 2.6556202608826744e-10 0 2.705620260882674e-10 0.00041 2.755620260882674e-10 0 2.659320680761243e-10 0 2.709320680761243e-10 0.00041 2.7593206807612427e-10 0 2.6728537619829637e-10 0 2.7228537619829635e-10 0.00041 2.7728537619829634e-10 0 2.775873572648208e-10 0 2.825873572648208e-10 0.00041 2.8758735726482077e-10 0 2.853328394445528e-10 0 2.9033283944455277e-10 0.00041 2.9533283944455276e-10 0 3.0270962454495933e-10 0 3.077096245449593e-10 0.00041 3.127096245449593e-10 0 3.068463254033064e-10 0 3.1184632540330636e-10 0.00041 3.1684632540330635e-10 0 3.113284330367877e-10 0 3.1632843303678767e-10 0.00041 3.2132843303678765e-10 0 3.298493565665906e-10 0 3.348493565665906e-10 0.00041 3.398493565665906e-10 0 3.4710149266782073e-10 0 3.521014926678207e-10 0.00041 3.571014926678207e-10 0 3.503360854033267e-10 0 3.5533608540332667e-10 0.00041 3.6033608540332665e-10 0 3.524436996121096e-10 0 3.5744369961210957e-10 0.00041 3.6244369961210956e-10 0 3.646766392097994e-10 0 3.6967663920979936e-10 0.00041 3.7467663920979934e-10 0 3.700598812425032e-10 0 3.7505988124250317e-10 0.00041 3.8005988124250315e-10 0 3.786067321796768e-10 0 3.836067321796768e-10 0.00041 3.886067321796768e-10 0 3.8909395428237484e-10 0 3.9409395428237483e-10 0.00041 3.990939542823748e-10 0 4.0141566072135247e-10 0 4.0641566072135245e-10 0.00041 4.1141566072135243e-10 0 4.306973538544831e-10 0 4.356973538544831e-10 0.00041 4.4069735385448306e-10 0 4.322342414403645e-10 0 4.372342414403645e-10 0.00041 4.422342414403645e-10 0 4.468922905922227e-10 0 4.518922905922227e-10 0.00041 4.568922905922227e-10 0 4.581346658829152e-10 0 4.631346658829152e-10 0.00041 4.681346658829152e-10 0 4.771151700662107e-10 0 4.821151700662107e-10 0.00041 4.871151700662107e-10 0 4.831050898076728e-10 0 4.881050898076728e-10 0.00041 4.931050898076728e-10 0 4.877919364508718e-10 0 4.927919364508717e-10 0.00041 4.977919364508717e-10 0 4.959630096156474e-10 0 5.009630096156474e-10 0.00041 5.059630096156474e-10 0 4.986077023991868e-10 0 5.036077023991868e-10 0.00041 5.086077023991868e-10 0 5.06065927289239e-10 0 5.11065927289239e-10 0.00041 5.16065927289239e-10 0 5.071265478490253e-10 0 5.121265478490253e-10 0.00041 5.171265478490253e-10 0 5.235960217857286e-10 0 5.285960217857285e-10 0.00041 5.335960217857285e-10 0 5.463884034615215e-10 0 5.513884034615215e-10 0.00041 5.563884034615215e-10 0 5.519094282069006e-10 0 5.569094282069006e-10 0.00041 5.619094282069005e-10 0 5.835367377340053e-10 0 5.885367377340053e-10 0.00041 5.935367377340053e-10 0 5.846137640484927e-10 0 5.896137640484927e-10 0.00041 5.946137640484927e-10 0 5.874091919557479e-10 0 5.924091919557479e-10 0.00041 5.974091919557479e-10 0 5.903816787860721e-10 0 5.953816787860721e-10 0.00041 6.003816787860721e-10 0 5.980172481553577e-10 0 6.030172481553577e-10 0.00041 6.080172481553576e-10 0 6.07374700760351e-10 0 6.12374700760351e-10 0.00041 6.17374700760351e-10 0 6.127341288681853e-10 0 6.177341288681853e-10 0.00041 6.227341288681853e-10 0 6.139796692092079e-10 0 6.189796692092078e-10 0.00041 6.239796692092078e-10 0 6.339595827749054e-10 0 6.389595827749054e-10 0.00041 6.439595827749054e-10 0 6.389342219294889e-10 0 6.439342219294889e-10 0.00041 6.489342219294889e-10 0 6.400699210760943e-10 0 6.450699210760942e-10 0.00041 6.500699210760942e-10 0 6.477822853514718e-10 0 6.527822853514718e-10 0.00041 6.577822853514718e-10 0 )
X32 SYNAPSE 31 0 32
X33 CONFLU 26 0 0 0 33
X34 CONFLU 23 28 30 32 34
X35 NEURON 33 34 35
IB36 8 0 pwl(0 0 5p 118.443u)
X37 SYNAPSE 8 0 37
IB38 12 0 pwl(0 0 5p 122.278u)
X39 SYNAPSE 12 0 39
IB40 16 0 pwl(0 0 5p 119.082u)
X41 SYNAPSE 0 16 41
IB43 20 0 pwl(0 0 5p 118.443u)
X44 SYNAPSE 20 0 44
IB45 45 0 pwl(0 0 5p 119.314u)
VIN45 45 0 pwl(0 0 1.7993190396890958e-12 0 6.7993190396890955e-12 0.00041 1.1799319039689095e-11 0 1.1995290054347743e-11 0 1.6995290054347742e-11 0.00041 2.199529005434774e-11 0 1.2193356680238297e-11 0 1.7193356680238296e-11 0.00041 2.2193356680238295e-11 0 1.2216049947050578e-11 0 1.7216049947050577e-11 0.00041 2.2216049947050576e-11 0 1.771947867344106e-11 0 2.271947867344106e-11 0.00041 2.7719478673441058e-11 0 3.401888302002491e-11 0 3.901888302002491e-11 0.00041 4.4018883020024913e-11 0 4.0754712546697226e-11 0 4.575471254669723e-11 0.00041 5.075471254669723e-11 0 4.8307726124951136e-11 0 5.330772612495114e-11 0.00041 5.830772612495113e-11 0 7.64755859157084e-11 0 8.147558591570839e-11 0.00041 8.647558591570839e-11 0 1.370531167201341e-10 0 1.4205311672013412e-10 0.00041 1.4705311672013412e-10 0 1.6991739929907154e-10 0 1.7491739929907155e-10 0.00041 1.7991739929907156e-10 0 1.6993027680241977e-10 0 1.7493027680241978e-10 0.00041 1.7993027680241979e-10 0 1.9262122344508884e-10 0 1.9762122344508885e-10 0.00041 2.0262122344508886e-10 0 1.9334620029428777e-10 0 1.9834620029428777e-10 0.00041 2.0334620029428778e-10 0 2.0404020331596094e-10 0 2.0904020331596095e-10 0.00041 2.1404020331596096e-10 0 2.125295336114063e-10 0 2.1752953361140632e-10 0.00041 2.2252953361140632e-10 0 2.440286201387913e-10 0 2.4902862013879126e-10 0.00041 2.5402862013879124e-10 0 2.4756872056072375e-10 0 2.5256872056072374e-10 0.00041 2.575687205607237e-10 0 2.506398319570072e-10 0 2.556398319570072e-10 0.00041 2.606398319570072e-10 0 2.6556202608826744e-10 0 2.705620260882674e-10 0.00041 2.755620260882674e-10 0 2.659320680761243e-10 0 2.709320680761243e-10 0.00041 2.7593206807612427e-10 0 2.6728537619829637e-10 0 2.7228537619829635e-10 0.00041 2.7728537619829634e-10 0 2.775873572648208e-10 0 2.825873572648208e-10 0.00041 2.8758735726482077e-10 0 2.853328394445528e-10 0 2.9033283944455277e-10 0.00041 2.9533283944455276e-10 0 3.0270962454495933e-10 0 3.077096245449593e-10 0.00041 3.127096245449593e-10 0 3.068463254033064e-10 0 3.1184632540330636e-10 0.00041 3.1684632540330635e-10 0 3.113284330367877e-10 0 3.1632843303678767e-10 0.00041 3.2132843303678765e-10 0 3.298493565665906e-10 0 3.348493565665906e-10 0.00041 3.398493565665906e-10 0 3.4710149266782073e-10 0 3.521014926678207e-10 0.00041 3.571014926678207e-10 0 3.503360854033267e-10 0 3.5533608540332667e-10 0.00041 3.6033608540332665e-10 0 3.524436996121096e-10 0 3.5744369961210957e-10 0.00041 3.6244369961210956e-10 0 3.646766392097994e-10 0 3.6967663920979936e-10 0.00041 3.7467663920979934e-10 0 3.700598812425032e-10 0 3.7505988124250317e-10 0.00041 3.8005988124250315e-10 0 3.786067321796768e-10 0 3.836067321796768e-10 0.00041 3.886067321796768e-10 0 3.8909395428237484e-10 0 3.9409395428237483e-10 0.00041 3.990939542823748e-10 0 4.0141566072135247e-10 0 4.0641566072135245e-10 0.00041 4.1141566072135243e-10 0 4.306973538544831e-10 0 4.356973538544831e-10 0.00041 4.4069735385448306e-10 0 4.322342414403645e-10 0 4.372342414403645e-10 0.00041 4.422342414403645e-10 0 4.468922905922227e-10 0 4.518922905922227e-10 0.00041 4.568922905922227e-10 0 4.581346658829152e-10 0 4.631346658829152e-10 0.00041 4.681346658829152e-10 0 4.771151700662107e-10 0 4.821151700662107e-10 0.00041 4.871151700662107e-10 0 4.831050898076728e-10 0 4.881050898076728e-10 0.00041 4.931050898076728e-10 0 4.877919364508718e-10 0 4.927919364508717e-10 0.00041 4.977919364508717e-10 0 4.959630096156474e-10 0 5.009630096156474e-10 0.00041 5.059630096156474e-10 0 4.986077023991868e-10 0 5.036077023991868e-10 0.00041 5.086077023991868e-10 0 5.06065927289239e-10 0 5.11065927289239e-10 0.00041 5.16065927289239e-10 0 5.071265478490253e-10 0 5.121265478490253e-10 0.00041 5.171265478490253e-10 0 5.235960217857286e-10 0 5.285960217857285e-10 0.00041 5.335960217857285e-10 0 5.463884034615215e-10 0 5.513884034615215e-10 0.00041 5.563884034615215e-10 0 5.519094282069006e-10 0 5.569094282069006e-10 0.00041 5.619094282069005e-10 0 5.835367377340053e-10 0 5.885367377340053e-10 0.00041 5.935367377340053e-10 0 5.846137640484927e-10 0 5.896137640484927e-10 0.00041 5.946137640484927e-10 0 5.874091919557479e-10 0 5.924091919557479e-10 0.00041 5.974091919557479e-10 0 5.903816787860721e-10 0 5.953816787860721e-10 0.00041 6.003816787860721e-10 0 5.980172481553577e-10 0 6.030172481553577e-10 0.00041 6.080172481553576e-10 0 6.07374700760351e-10 0 6.12374700760351e-10 0.00041 6.17374700760351e-10 0 6.127341288681853e-10 0 6.177341288681853e-10 0.00041 6.227341288681853e-10 0 6.139796692092079e-10 0 6.189796692092078e-10 0.00041 6.239796692092078e-10 0 6.339595827749054e-10 0 6.389595827749054e-10 0.00041 6.439595827749054e-10 0 6.389342219294889e-10 0 6.439342219294889e-10 0.00041 6.489342219294889e-10 0 6.400699210760943e-10 0 6.450699210760942e-10 0.00041 6.500699210760942e-10 0 6.477822853514718e-10 0 6.527822853514718e-10 0.00041 6.577822853514718e-10 0 )
X46 SYNAPSE 45 0 46
X47 CONFLU 42 0 0 0 47
X48 CONFLU 37 39 44 46 48
X49 NEURON 47 48 49
IB50 9 0 pwl(0 0 5p 116.753u)
X51 SYNAPSE 0 9 51
IB53 13 0 pwl(0 0 5p 118.378u)
X54 SYNAPSE 13 0 54
IB55 17 0 pwl(0 0 5p 121.273u)
X56 SYNAPSE 0 17 56
IB58 21 0 pwl(0 0 5p 134.829u)
X59 SYNAPSE 0 21 59
IB61 61 0 pwl(0 0 5p 117.972u)
VIN61 61 0 pwl(0 0 1.7993190396890958e-12 0 6.7993190396890955e-12 0.00041 1.1799319039689095e-11 0 1.1995290054347743e-11 0 1.6995290054347742e-11 0.00041 2.199529005434774e-11 0 1.2193356680238297e-11 0 1.7193356680238296e-11 0.00041 2.2193356680238295e-11 0 1.2216049947050578e-11 0 1.7216049947050577e-11 0.00041 2.2216049947050576e-11 0 1.771947867344106e-11 0 2.271947867344106e-11 0.00041 2.7719478673441058e-11 0 3.401888302002491e-11 0 3.901888302002491e-11 0.00041 4.4018883020024913e-11 0 4.0754712546697226e-11 0 4.575471254669723e-11 0.00041 5.075471254669723e-11 0 4.8307726124951136e-11 0 5.330772612495114e-11 0.00041 5.830772612495113e-11 0 7.64755859157084e-11 0 8.147558591570839e-11 0.00041 8.647558591570839e-11 0 1.370531167201341e-10 0 1.4205311672013412e-10 0.00041 1.4705311672013412e-10 0 1.6991739929907154e-10 0 1.7491739929907155e-10 0.00041 1.7991739929907156e-10 0 1.6993027680241977e-10 0 1.7493027680241978e-10 0.00041 1.7993027680241979e-10 0 1.9262122344508884e-10 0 1.9762122344508885e-10 0.00041 2.0262122344508886e-10 0 1.9334620029428777e-10 0 1.9834620029428777e-10 0.00041 2.0334620029428778e-10 0 2.0404020331596094e-10 0 2.0904020331596095e-10 0.00041 2.1404020331596096e-10 0 2.125295336114063e-10 0 2.1752953361140632e-10 0.00041 2.2252953361140632e-10 0 2.440286201387913e-10 0 2.4902862013879126e-10 0.00041 2.5402862013879124e-10 0 2.4756872056072375e-10 0 2.5256872056072374e-10 0.00041 2.575687205607237e-10 0 2.506398319570072e-10 0 2.556398319570072e-10 0.00041 2.606398319570072e-10 0 2.6556202608826744e-10 0 2.705620260882674e-10 0.00041 2.755620260882674e-10 0 2.659320680761243e-10 0 2.709320680761243e-10 0.00041 2.7593206807612427e-10 0 2.6728537619829637e-10 0 2.7228537619829635e-10 0.00041 2.7728537619829634e-10 0 2.775873572648208e-10 0 2.825873572648208e-10 0.00041 2.8758735726482077e-10 0 2.853328394445528e-10 0 2.9033283944455277e-10 0.00041 2.9533283944455276e-10 0 3.0270962454495933e-10 0 3.077096245449593e-10 0.00041 3.127096245449593e-10 0 3.068463254033064e-10 0 3.1184632540330636e-10 0.00041 3.1684632540330635e-10 0 3.113284330367877e-10 0 3.1632843303678767e-10 0.00041 3.2132843303678765e-10 0 3.298493565665906e-10 0 3.348493565665906e-10 0.00041 3.398493565665906e-10 0 3.4710149266782073e-10 0 3.521014926678207e-10 0.00041 3.571014926678207e-10 0 3.503360854033267e-10 0 3.5533608540332667e-10 0.00041 3.6033608540332665e-10 0 3.524436996121096e-10 0 3.5744369961210957e-10 0.00041 3.6244369961210956e-10 0 3.646766392097994e-10 0 3.6967663920979936e-10 0.00041 3.7467663920979934e-10 0 3.700598812425032e-10 0 3.7505988124250317e-10 0.00041 3.8005988124250315e-10 0 3.786067321796768e-10 0 3.836067321796768e-10 0.00041 3.886067321796768e-10 0 3.8909395428237484e-10 0 3.9409395428237483e-10 0.00041 3.990939542823748e-10 0 4.0141566072135247e-10 0 4.0641566072135245e-10 0.00041 4.1141566072135243e-10 0 4.306973538544831e-10 0 4.356973538544831e-10 0.00041 4.4069735385448306e-10 0 4.322342414403645e-10 0 4.372342414403645e-10 0.00041 4.422342414403645e-10 0 4.468922905922227e-10 0 4.518922905922227e-10 0.00041 4.568922905922227e-10 0 4.581346658829152e-10 0 4.631346658829152e-10 0.00041 4.681346658829152e-10 0 4.771151700662107e-10 0 4.821151700662107e-10 0.00041 4.871151700662107e-10 0 4.831050898076728e-10 0 4.881050898076728e-10 0.00041 4.931050898076728e-10 0 4.877919364508718e-10 0 4.927919364508717e-10 0.00041 4.977919364508717e-10 0 4.959630096156474e-10 0 5.009630096156474e-10 0.00041 5.059630096156474e-10 0 4.986077023991868e-10 0 5.036077023991868e-10 0.00041 5.086077023991868e-10 0 5.06065927289239e-10 0 5.11065927289239e-10 0.00041 5.16065927289239e-10 0 5.071265478490253e-10 0 5.121265478490253e-10 0.00041 5.171265478490253e-10 0 5.235960217857286e-10 0 5.285960217857285e-10 0.00041 5.335960217857285e-10 0 5.463884034615215e-10 0 5.513884034615215e-10 0.00041 5.563884034615215e-10 0 5.519094282069006e-10 0 5.569094282069006e-10 0.00041 5.619094282069005e-10 0 5.835367377340053e-10 0 5.885367377340053e-10 0.00041 5.935367377340053e-10 0 5.846137640484927e-10 0 5.896137640484927e-10 0.00041 5.946137640484927e-10 0 5.874091919557479e-10 0 5.924091919557479e-10 0.00041 5.974091919557479e-10 0 5.903816787860721e-10 0 5.953816787860721e-10 0.00041 6.003816787860721e-10 0 5.980172481553577e-10 0 6.030172481553577e-10 0.00041 6.080172481553576e-10 0 6.07374700760351e-10 0 6.12374700760351e-10 0.00041 6.17374700760351e-10 0 6.127341288681853e-10 0 6.177341288681853e-10 0.00041 6.227341288681853e-10 0 6.139796692092079e-10 0 6.189796692092078e-10 0.00041 6.239796692092078e-10 0 6.339595827749054e-10 0 6.389595827749054e-10 0.00041 6.439595827749054e-10 0 6.389342219294889e-10 0 6.439342219294889e-10 0.00041 6.489342219294889e-10 0 6.400699210760943e-10 0 6.450699210760942e-10 0.00041 6.500699210760942e-10 0 6.477822853514718e-10 0 6.527822853514718e-10 0.00041 6.577822853514718e-10 0 )
X62 SYNAPSE 0 61 62
X63 CONFLU 52 57 60 62 63
X64 CONFLU 54 0 0 0 64
X65 NEURON 63 64 65
.temp 4.2
    .model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
    .tran 0.008 220p 0 0.008p
    .print PHASE 35 0
.print PHASE 49 0
.print PHASE 65 0
.end