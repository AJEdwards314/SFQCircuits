.subckt DCSFQ 2 17
B01        5          3          jj1     area=1.32
B02        5          6          jj1     area=1
B03        9          10         jj1     area=1.5
B04        13         14         jj1     area=1.96
B05        15         16         jj1     area=1.96
IB01       0          8          pwl(0 0 5p 162.5u)
IB02       0          12         pwl(0 0 5p 260u)
L01        2          1          0.848p
L02        0          1          7.712p
L03        1          3          1.778p
L04        5          7          0.543p
L05        7          9          3.149p
L06        9          11         1.323p
L07        11         13         1.095p
L08        13         15         2.951p
L09        15         17         1.63p
LP01       0          6          0.398p
LP02       0          10         0.211p
LP03       0          14         0.276p
LP04       0          16         0.224p
LPR01      7          8          0.915p
LPR02      11         12         0.307p
LRB01      4          5          1p
LRB02      18         6          1p
LRB03      19         10         1p
LRB04      20         14         1p
LRB05      21         16         1p
RB01       3          4          8.56
RB02       18         5          11.30
RB03       19         9          7.53
RB04       20         13         5.77
RB05       21         15         5.77
.model jj1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.ends DCSFQ

.subckt CONFLU 1 2 3 4 14
B01 5 0 jmitll
B02 5 9 jmitll area=1.5
B03 6 0 jmitll
B04 6 10 jmitll area=1.5
B05 7 0 jmitll
B06 7 11 jmitll area=1.5
B07 8 0 jmitll
B08 8 12 jmitll area=1.5
B0L 14 0 jmitll
L01 1 5 0.5p
L02 2 6 0.5p
L03 3 7 0.5p
L04 4 8 0.5p
L05 9 13 0.5p
L06 10 13 0.5p
L07 11 13 0.5p
L08 12 13 0.5p
LC1 13 14 2p
I01 0 13 pwl(0 0 5p 800u)
.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.ends CONFLU

.subckt NEURON 11 5 4
B01        0          11         jmitll
B02        0          4          jmitll
B03        0          5          jmitll
IB0        0          11         pwl(0 0 5p 0u)
L02        11         2          5p
L03        5          6          5p
L04        3          4          5p
K01        L04        L03        0.6
R01        2          3          0.5
R02        3          0          0.075
R03        6          0          0.2
.ends NEURON

.subckt SYNAPSE 1 6 7
B01        7          1          jmitll
B02        0          7          jmitll
L01        7          9          0.1p
L02        6          7          0.1p
.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
.ends SYNAPSE

.subckt SPLITTER 1 3 4
* Splitting Circuit w/ Output Buffers

# Junctions
B01	2	0	 jmitll
B02	4	0	 jmitll
B03	5	0	 jmitll
B04	6	0	 jmitll
B05	7	0	 jmitll
B06	6	8	 jmitll2
B07	7	9	 jmitll2

# Inductors
L01	1	2	0.5p
L02	2	3	0.5p
L03	3	5	0.5p
L04	3	4	0.5p
L05	5	7	0.5p
L06	4	6	0.5p
L07	9	11	0.5p
L08	8	10	0.5p

# Bias Currents
I01	3	0	 pwl(0 0 5p 250u)
I02	9	0	 pwl(0 0 5p 175u)
I03	8	0	 pwl(0 0 5p 175u)

# Resistors
R0L1    11  0   1
R0L2    10  0   1
R0L     3   0   1

.model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.2mA)
.model jmitll2 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.1mA)
.ends SPLITTER
VIN1 1 0 pwl(0 0 5.298467839300459e-12 0 1.5298467839300458e-11 0.00021 2.5298467839300456e-11 0 2.8239402622282406e-11 0 3.8239402622282403e-11 0.00021 4.82394026222824e-11 0 4.823940262228241e-11 0 5.82394026222824e-11 0.00021 6.823940262228241e-11 0 6.82394026222824e-11 0 7.82394026222824e-11 0.00021 8.82394026222824e-11 0 8.82394026222824e-11 0 9.823940262228241e-11 0.00021 1.0823940262228241e-10 0 1.0823940262228239e-10 0 1.182394026222824e-10 0.00021 1.2823940262228238e-10 0 1.2823940262228238e-10 0 1.3823940262228237e-10 0.00021 1.4823940262228237e-10 0 1.4823940262228237e-10 0 1.5823940262228236e-10 0.00021 1.6823940262228235e-10 0 1.733200683103438e-10 0 1.833200683103438e-10 0.00021 1.933200683103438e-10 0 3.096195126203016e-10 0 3.196195126203016e-10 0.00021 3.2961951262030163e-10 0 3.835641484229108e-10 0 3.935641484229108e-10 0.00021 4.035641484229108e-10 0 4.0356414842291076e-10 0 4.135641484229108e-10 0.00021 4.235641484229108e-10 0 4.346477527514497e-10 0 4.446477527514497e-10 0.00021 4.546477527514497e-10 0 4.5464775275144966e-10 0 4.646477527514497e-10 0.00021 4.746477527514496e-10 0 4.746477527514498e-10 0 4.846477527514497e-10 0.00021 4.946477527514497e-10 0 4.946477527514498e-10 0 5.046477527514498e-10 0.00021 5.146477527514497e-10 0 )
VIN2 2 0 pwl(0 0 2.3996595198445482e-11 0 3.399659519844548e-11 0.00021 4.399659519844548e-11 0 7.497645027173871e-11 0 8.497645027173871e-11 0.00021 9.497645027173872e-11 0 9.49764502717387e-11 0 1.0497645027173871e-10 0.00021 1.1497645027173871e-10 0 1.149764502717387e-10 0 1.249764502717387e-10 0.00021 1.349764502717387e-10 0 1.3497645027173872e-10 0 1.449764502717387e-10 0.00021 1.549764502717387e-10 0 1.8509441510012458e-10 0 1.9509441510012457e-10 0.00021 2.0509441510012456e-10 0 2.1877356273348619e-10 0 2.2877356273348618e-10 0.00021 2.387735627334862e-10 0 2.5653863062475574e-10 0 2.6653863062475575e-10 0.00021 2.7653863062475577e-10 0 3.9737792957854203e-10 0 4.0737792957854204e-10 0.00021 4.1737792957854206e-10 0 )
VIN3 3 0 pwl(0 0 -1.6765138868488735e-13 0 9.832348611315112e-12 0.00021 1.983234861131511e-11 0 1.9832348611315116e-11 0 2.9832348611315114e-11 0.00021 3.983234861131511e-11 0 3.983234861131511e-11 0 4.983234861131511e-11 0.00021 5.983234861131511e-11 0 5.98323486113151e-11 0 6.98323486113151e-11 0.00021 7.983234861131511e-11 0 7.98323486113151e-11 0 8.98323486113151e-11 0.00021 9.98323486113151e-11 0 9.983234861131509e-11 0 1.098323486113151e-10 0.00021 1.198323486113151e-10 0 1.1983234861131511e-10 0 1.298323486113151e-10 0.00021 1.398323486113151e-10 0 1.398323486113151e-10 0 1.498323486113151e-10 0.00021 1.5983234861131508e-10 0 1.5983234861131508e-10 0 1.6983234861131507e-10 0.00021 1.7983234861131506e-10 0 1.9541994819823317e-10 0 2.0541994819823316e-10 0.00021 2.1541994819823315e-10 0 2.4294427839816715e-10 0 2.5294427839816717e-10 0.00021 2.629442783981672e-10 0 2.6294427839816714e-10 0 2.7294427839816715e-10 0.00021 2.8294427839816717e-10 0 2.829442783981671e-10 0 2.9294427839816714e-10 0.00021 3.0294427839816715e-10 0 3.029442783981671e-10 0 3.129442783981671e-10 0.00021 3.2294427839816714e-10 0 3.229442783981671e-10 0 3.329442783981671e-10 0.00021 3.429442783981671e-10 0 3.4294427839816707e-10 0 3.529442783981671e-10 0.00021 3.629442783981671e-10 0 3.6294427839816705e-10 0 3.7294427839816707e-10 0.00021 3.829442783981671e-10 0 3.8294427839816703e-10 0 3.9294427839816705e-10 0.00021 4.0294427839816707e-10 0 4.02944278398167e-10 0 4.1294427839816703e-10 0.00021 4.2294427839816705e-10 0 4.22944278398167e-10 0 4.32944278398167e-10 0.00021 4.4294427839816703e-10 0 4.42944278398167e-10 0 4.52944278398167e-10 0.00021 4.62944278398167e-10 0 4.6294427839816696e-10 0 4.72944278398167e-10 0.00021 4.829442783981669e-10 0 4.82944278398167e-10 0 4.92944278398167e-10 0.00021 5.02944278398167e-10 0 5.029442783981671e-10 0 5.12944278398167e-10 0.00021 5.22944278398167e-10 0 5.229442783981671e-10 0 5.329442783981671e-10 0.00021 5.42944278398167e-10 0 5.429442783981672e-10 0 5.529442783981671e-10 0.00021 5.629442783981671e-10 0 5.629442783981672e-10 0 5.729442783981672e-10 0.00021 5.829442783981671e-10 0 5.829442783981672e-10 0 5.929442783981672e-10 0.00021 6.029442783981672e-10 0 )
VIN4 4 0 pwl(0 0 -7.282013095148655e-13 0 9.271798690485134e-12 0.00021 1.9271798690485132e-11 0 1.9271798690485138e-11 0 2.9271798690485136e-11 0.00021 3.9271798690485134e-11 0 3.9271798690485134e-11 0 4.927179869048513e-11 0.00021 5.927179869048514e-11 0 5.927179869048512e-11 0 6.927179869048513e-11 0.00021 7.927179869048513e-11 0 7.927179869048512e-11 0 8.927179869048512e-11 0.00021 9.927179869048513e-11 0 9.927179869048513e-11 0 1.0927179869048513e-10 0.00021 1.1927179869048512e-10 0 1.1927179869048512e-10 0 1.2927179869048511e-10 0.00021 1.392717986904851e-10 0 1.392717986904851e-10 0 1.492717986904851e-10 0.00021 1.592717986904851e-10 0 1.592717986904851e-10 0 1.6927179869048508e-10 0.00021 1.7927179869048507e-10 0 1.837087955274557e-10 0 1.937087955274557e-10 0.00021 2.037087955274557e-10 0 2.2852372631691587e-10 0 2.3852372631691586e-10 0.00021 2.485237263169159e-10 0 2.485237263169158e-10 0 2.5852372631691584e-10 0.00021 2.6852372631691586e-10 0 2.685237263169158e-10 0 2.785237263169158e-10 0.00021 2.8852372631691584e-10 0 2.885237263169158e-10 0 2.985237263169158e-10 0.00021 3.085237263169158e-10 0 3.0852372631691577e-10 0 3.185237263169158e-10 0.00021 3.285237263169158e-10 0 3.2852372631691576e-10 0 3.3852372631691577e-10 0.00021 3.485237263169158e-10 0 3.4852372631691574e-10 0 3.5852372631691576e-10 0.00021 3.6852372631691577e-10 0 3.685237263169157e-10 0 3.7852372631691574e-10 0.00021 3.8852372631691576e-10 0 3.885237263169157e-10 0 3.985237263169157e-10 0.00021 4.0852372631691574e-10 0 4.085237263169157e-10 0 4.185237263169157e-10 0.00021 4.285237263169157e-10 0 4.2852372631691567e-10 0 4.385237263169157e-10 0.00021 4.485237263169157e-10 0 4.4852372631691565e-10 0 4.5852372631691567e-10 0.00021 4.685237263169157e-10 0 4.685237263169157e-10 0 4.785237263169157e-10 0.00021 4.885237263169156e-10 0 4.885237263169157e-10 0 4.985237263169157e-10 0.00021 5.085237263169157e-10 0 5.085237263169158e-10 0 5.185237263169157e-10 0.00021 5.285237263169157e-10 0 5.285237263169158e-10 0 5.385237263169158e-10 0.00021 5.485237263169157e-10 0 5.485237263169158e-10 0 5.585237263169158e-10 0.00021 5.685237263169158e-10 0 5.685237263169159e-10 0 5.785237263169158e-10 0.00021 5.885237263169158e-10 0 5.885237263169159e-10 0 5.985237263169159e-10 0.00021 6.085237263169158e-10 0 6.085237263169159e-10 0 6.185237263169159e-10 0.00021 6.285237263169159e-10 0 6.28523726316916e-10 0 6.385237263169159e-10 0.00021 6.485237263169159e-10 0 )
VIN5 5 0 pwl(0 0 -1.5008512003886294e-12 0 8.49914879961137e-12 0.00021 1.8499148799611368e-11 0 1.8499148799611368e-11 0 2.849914879961137e-11 0.00021 3.849914879961137e-11 0 3.849914879961137e-11 0 4.849914879961137e-11 0.00021 5.849914879961137e-11 0 5.849914879961136e-11 0 6.849914879961136e-11 0.00021 7.849914879961137e-11 0 7.849914879961135e-11 0 8.849914879961136e-11 0.00021 9.849914879961136e-11 0 9.849914879961136e-11 0 1.0849914879961137e-10 0.00021 1.1849914879961136e-10 0 1.1849914879961138e-10 0 1.2849914879961138e-10 0.00021 1.3849914879961137e-10 0 1.3849914879961137e-10 0 1.4849914879961136e-10 0.00021 1.5849914879961135e-10 0 1.5849914879961135e-10 0 1.6849914879961134e-10 0.00021 1.7849914879961133e-10 0 1.7849914879961136e-10 0 1.8849914879961135e-10 0.00021 1.9849914879961134e-10 0 2.0864674912383949e-10 0 2.1864674912383948e-10 0.00021 2.2864674912383947e-10 0 2.286467491238395e-10 0 2.386467491238395e-10 0.00021 2.486467491238395e-10 0 2.4864674912383945e-10 0 2.5864674912383947e-10 0.00021 2.686467491238395e-10 0 2.6864674912383943e-10 0 2.7864674912383945e-10 0.00021 2.8864674912383947e-10 0 2.886467491238394e-10 0 2.9864674912383943e-10 0.00021 3.0864674912383945e-10 0 3.086467491238394e-10 0 3.186467491238394e-10 0.00021 3.2864674912383943e-10 0 3.286467491238394e-10 0 3.386467491238394e-10 0.00021 3.486467491238394e-10 0 3.4864674912383936e-10 0 3.586467491238394e-10 0.00021 3.686467491238394e-10 0 3.6864674912383935e-10 0 3.7864674912383936e-10 0.00021 3.886467491238394e-10 0 3.8864674912383933e-10 0 3.9864674912383935e-10 0.00021 4.0864674912383936e-10 0 4.086467491238393e-10 0 4.1864674912383933e-10 0.00021 4.2864674912383935e-10 0 4.286467491238393e-10 0 4.386467491238393e-10 0.00021 4.4864674912383933e-10 0 4.486467491238393e-10 0 4.586467491238393e-10 0.00021 4.686467491238393e-10 0 4.686467491238394e-10 0 4.786467491238393e-10 0.00021 4.886467491238393e-10 0 4.886467491238394e-10 0 4.986467491238394e-10 0.00021 5.086467491238393e-10 0 5.086467491238394e-10 0 5.186467491238394e-10 0.00021 5.286467491238394e-10 0 5.286467491238395e-10 0 5.386467491238394e-10 0.00021 5.486467491238394e-10 0 5.486467491238395e-10 0 5.586467491238395e-10 0.00021 5.686467491238394e-10 0 5.686467491238395e-10 0 5.786467491238395e-10 0.00021 5.886467491238395e-10 0 5.886467491238396e-10 0 5.986467491238395e-10 0.00021 6.086467491238395e-10 0 6.086467491238396e-10 0 6.186467491238396e-10 0.00021 6.286467491238395e-10 0 6.286467491238396e-10 0 6.386467491238396e-10 0.00021 6.486467491238396e-10 0 6.486467491238397e-10 0 6.586467491238396e-10 0.00021 6.686467491238396e-10 0 6.686467491238397e-10 0 6.786467491238397e-10 0.00021 6.886467491238396e-10 0 6.886467491238397e-10 0 6.986467491238397e-10 0.00021 7.086467491238397e-10 0 )
X6 SPLITTER 1 6 7
X7 SPLITTER 7 8 9
X8 SPLITTER 2 10 11
X9 SPLITTER 11 12 13
X10 SPLITTER 3 14 15
X11 SPLITTER 15 16 17
X12 SPLITTER 4 18 19
X13 SPLITTER 19 20 21
IB22 22 0 pwl(0 0 5p 120.946u)
X23 SYNAPSE 6 22 23
IB24 24 0 pwl(0 0 5p 120.242u)
X25 SYNAPSE 10 24 25
IB27 27 0 pwl(0 0 5p 119.076u)
X28 SYNAPSE 14 27 28
IB29 29 0 pwl(0 0 5p 124.75u)
X30 SYNAPSE 18 29 30
IB31 31 0 pwl(0 0 5p 118.06u)
VIN32 32 0 pwl(0 0 -1.5008512003886294e-12 0 8.49914879961137e-12 0.00021 1.8499148799611368e-11 0 1.8499148799611368e-11 0 2.849914879961137e-11 0.00021 3.849914879961137e-11 0 3.849914879961137e-11 0 4.849914879961137e-11 0.00021 5.849914879961137e-11 0 5.849914879961136e-11 0 6.849914879961136e-11 0.00021 7.849914879961137e-11 0 7.849914879961135e-11 0 8.849914879961136e-11 0.00021 9.849914879961136e-11 0 9.849914879961136e-11 0 1.0849914879961137e-10 0.00021 1.1849914879961136e-10 0 1.1849914879961138e-10 0 1.2849914879961138e-10 0.00021 1.3849914879961137e-10 0 1.3849914879961137e-10 0 1.4849914879961136e-10 0.00021 1.5849914879961135e-10 0 1.5849914879961135e-10 0 1.6849914879961134e-10 0.00021 1.7849914879961133e-10 0 1.7849914879961136e-10 0 1.8849914879961135e-10 0.00021 1.9849914879961134e-10 0 2.0864674912383949e-10 0 2.1864674912383948e-10 0.00021 2.2864674912383947e-10 0 2.286467491238395e-10 0 2.386467491238395e-10 0.00021 2.486467491238395e-10 0 2.4864674912383945e-10 0 2.5864674912383947e-10 0.00021 2.686467491238395e-10 0 2.6864674912383943e-10 0 2.7864674912383945e-10 0.00021 2.8864674912383947e-10 0 2.886467491238394e-10 0 2.9864674912383943e-10 0.00021 3.0864674912383945e-10 0 3.086467491238394e-10 0 3.186467491238394e-10 0.00021 3.2864674912383943e-10 0 3.286467491238394e-10 0 3.386467491238394e-10 0.00021 3.486467491238394e-10 0 3.4864674912383936e-10 0 3.586467491238394e-10 0.00021 3.686467491238394e-10 0 3.6864674912383935e-10 0 3.7864674912383936e-10 0.00021 3.886467491238394e-10 0 3.8864674912383933e-10 0 3.9864674912383935e-10 0.00021 4.0864674912383936e-10 0 4.086467491238393e-10 0 4.1864674912383933e-10 0.00021 4.2864674912383935e-10 0 4.286467491238393e-10 0 4.386467491238393e-10 0.00021 4.4864674912383933e-10 0 4.486467491238393e-10 0 4.586467491238393e-10 0.00021 4.686467491238393e-10 0 4.686467491238394e-10 0 4.786467491238393e-10 0.00021 4.886467491238393e-10 0 4.886467491238394e-10 0 4.986467491238394e-10 0.00021 5.086467491238393e-10 0 5.086467491238394e-10 0 5.186467491238394e-10 0.00021 5.286467491238394e-10 0 5.286467491238395e-10 0 5.386467491238394e-10 0.00021 5.486467491238394e-10 0 5.486467491238395e-10 0 5.586467491238395e-10 0.00021 5.686467491238394e-10 0 5.686467491238395e-10 0 5.786467491238395e-10 0.00021 5.886467491238395e-10 0 5.886467491238396e-10 0 5.986467491238395e-10 0.00021 6.086467491238395e-10 0 6.086467491238396e-10 0 6.186467491238396e-10 0.00021 6.286467491238395e-10 0 6.286467491238396e-10 0 6.386467491238396e-10 0.00021 6.486467491238396e-10 0 6.486467491238397e-10 0 6.586467491238396e-10 0.00021 6.686467491238396e-10 0 6.686467491238397e-10 0 6.786467491238397e-10 0.00021 6.886467491238396e-10 0 6.886467491238397e-10 0 6.986467491238397e-10 0.00021 7.086467491238397e-10 0 )
X33 SYNAPSE 32 31 33
X35 CONFLU 23 28 30 33 35
X34 CONFLU 26 0 0 0 34
X36 NEURON 34 35 36
IB37 37 0 pwl(0 0 5p 118.098u)
X38 SYNAPSE 8 37 38
IB40 40 0 pwl(0 0 5p 122.37u)
X41 SYNAPSE 12 40 41
IB42 42 0 pwl(0 0 5p 118.679u)
X43 SYNAPSE 16 42 43
IB45 45 0 pwl(0 0 5p 119.513u)
X46 SYNAPSE 20 45 46
IB47 47 0 pwl(0 0 5p 119.364u)
VIN48 48 0 pwl(0 0 -1.5008512003886294e-12 0 8.49914879961137e-12 0.00021 1.8499148799611368e-11 0 1.8499148799611368e-11 0 2.849914879961137e-11 0.00021 3.849914879961137e-11 0 3.849914879961137e-11 0 4.849914879961137e-11 0.00021 5.849914879961137e-11 0 5.849914879961136e-11 0 6.849914879961136e-11 0.00021 7.849914879961137e-11 0 7.849914879961135e-11 0 8.849914879961136e-11 0.00021 9.849914879961136e-11 0 9.849914879961136e-11 0 1.0849914879961137e-10 0.00021 1.1849914879961136e-10 0 1.1849914879961138e-10 0 1.2849914879961138e-10 0.00021 1.3849914879961137e-10 0 1.3849914879961137e-10 0 1.4849914879961136e-10 0.00021 1.5849914879961135e-10 0 1.5849914879961135e-10 0 1.6849914879961134e-10 0.00021 1.7849914879961133e-10 0 1.7849914879961136e-10 0 1.8849914879961135e-10 0.00021 1.9849914879961134e-10 0 2.0864674912383949e-10 0 2.1864674912383948e-10 0.00021 2.2864674912383947e-10 0 2.286467491238395e-10 0 2.386467491238395e-10 0.00021 2.486467491238395e-10 0 2.4864674912383945e-10 0 2.5864674912383947e-10 0.00021 2.686467491238395e-10 0 2.6864674912383943e-10 0 2.7864674912383945e-10 0.00021 2.8864674912383947e-10 0 2.886467491238394e-10 0 2.9864674912383943e-10 0.00021 3.0864674912383945e-10 0 3.086467491238394e-10 0 3.186467491238394e-10 0.00021 3.2864674912383943e-10 0 3.286467491238394e-10 0 3.386467491238394e-10 0.00021 3.486467491238394e-10 0 3.4864674912383936e-10 0 3.586467491238394e-10 0.00021 3.686467491238394e-10 0 3.6864674912383935e-10 0 3.7864674912383936e-10 0.00021 3.886467491238394e-10 0 3.8864674912383933e-10 0 3.9864674912383935e-10 0.00021 4.0864674912383936e-10 0 4.086467491238393e-10 0 4.1864674912383933e-10 0.00021 4.2864674912383935e-10 0 4.286467491238393e-10 0 4.386467491238393e-10 0.00021 4.4864674912383933e-10 0 4.486467491238393e-10 0 4.586467491238393e-10 0.00021 4.686467491238393e-10 0 4.686467491238394e-10 0 4.786467491238393e-10 0.00021 4.886467491238393e-10 0 4.886467491238394e-10 0 4.986467491238394e-10 0.00021 5.086467491238393e-10 0 5.086467491238394e-10 0 5.186467491238394e-10 0.00021 5.286467491238394e-10 0 5.286467491238395e-10 0 5.386467491238394e-10 0.00021 5.486467491238394e-10 0 5.486467491238395e-10 0 5.586467491238395e-10 0.00021 5.686467491238394e-10 0 5.686467491238395e-10 0 5.786467491238395e-10 0.00021 5.886467491238395e-10 0 5.886467491238396e-10 0 5.986467491238395e-10 0.00021 6.086467491238395e-10 0 6.086467491238396e-10 0 6.186467491238396e-10 0.00021 6.286467491238395e-10 0 6.286467491238396e-10 0 6.386467491238396e-10 0.00021 6.486467491238396e-10 0 6.486467491238397e-10 0 6.586467491238396e-10 0.00021 6.686467491238396e-10 0 6.686467491238397e-10 0 6.786467491238397e-10 0.00021 6.886467491238396e-10 0 6.886467491238397e-10 0 6.986467491238397e-10 0.00021 7.086467491238397e-10 0 )
X49 SYNAPSE 48 47 49
X51 CONFLU 41 46 49 0 51
X50 CONFLU 39 44 0 0 50
X52 NEURON 50 51 52
IB53 53 0 pwl(0 0 5p 118.112u)
X54 SYNAPSE 9 53 54
IB56 56 0 pwl(0 0 5p 118.741u)
X57 SYNAPSE 13 56 57
IB58 58 0 pwl(0 0 5p 120.624u)
X59 SYNAPSE 17 58 59
IB61 61 0 pwl(0 0 5p 125.379u)
X62 SYNAPSE 21 61 62
IB64 64 0 pwl(0 0 5p 118.095u)
VIN65 65 0 pwl(0 0 -1.5008512003886294e-12 0 8.49914879961137e-12 0.00021 1.8499148799611368e-11 0 1.8499148799611368e-11 0 2.849914879961137e-11 0.00021 3.849914879961137e-11 0 3.849914879961137e-11 0 4.849914879961137e-11 0.00021 5.849914879961137e-11 0 5.849914879961136e-11 0 6.849914879961136e-11 0.00021 7.849914879961137e-11 0 7.849914879961135e-11 0 8.849914879961136e-11 0.00021 9.849914879961136e-11 0 9.849914879961136e-11 0 1.0849914879961137e-10 0.00021 1.1849914879961136e-10 0 1.1849914879961138e-10 0 1.2849914879961138e-10 0.00021 1.3849914879961137e-10 0 1.3849914879961137e-10 0 1.4849914879961136e-10 0.00021 1.5849914879961135e-10 0 1.5849914879961135e-10 0 1.6849914879961134e-10 0.00021 1.7849914879961133e-10 0 1.7849914879961136e-10 0 1.8849914879961135e-10 0.00021 1.9849914879961134e-10 0 2.0864674912383949e-10 0 2.1864674912383948e-10 0.00021 2.2864674912383947e-10 0 2.286467491238395e-10 0 2.386467491238395e-10 0.00021 2.486467491238395e-10 0 2.4864674912383945e-10 0 2.5864674912383947e-10 0.00021 2.686467491238395e-10 0 2.6864674912383943e-10 0 2.7864674912383945e-10 0.00021 2.8864674912383947e-10 0 2.886467491238394e-10 0 2.9864674912383943e-10 0.00021 3.0864674912383945e-10 0 3.086467491238394e-10 0 3.186467491238394e-10 0.00021 3.2864674912383943e-10 0 3.286467491238394e-10 0 3.386467491238394e-10 0.00021 3.486467491238394e-10 0 3.4864674912383936e-10 0 3.586467491238394e-10 0.00021 3.686467491238394e-10 0 3.6864674912383935e-10 0 3.7864674912383936e-10 0.00021 3.886467491238394e-10 0 3.8864674912383933e-10 0 3.9864674912383935e-10 0.00021 4.0864674912383936e-10 0 4.086467491238393e-10 0 4.1864674912383933e-10 0.00021 4.2864674912383935e-10 0 4.286467491238393e-10 0 4.386467491238393e-10 0.00021 4.4864674912383933e-10 0 4.486467491238393e-10 0 4.586467491238393e-10 0.00021 4.686467491238393e-10 0 4.686467491238394e-10 0 4.786467491238393e-10 0.00021 4.886467491238393e-10 0 4.886467491238394e-10 0 4.986467491238394e-10 0.00021 5.086467491238393e-10 0 5.086467491238394e-10 0 5.186467491238394e-10 0.00021 5.286467491238394e-10 0 5.286467491238395e-10 0 5.386467491238394e-10 0.00021 5.486467491238394e-10 0 5.486467491238395e-10 0 5.586467491238395e-10 0.00021 5.686467491238394e-10 0 5.686467491238395e-10 0 5.786467491238395e-10 0.00021 5.886467491238395e-10 0 5.886467491238396e-10 0 5.986467491238395e-10 0.00021 6.086467491238395e-10 0 6.086467491238396e-10 0 6.186467491238396e-10 0.00021 6.286467491238395e-10 0 6.286467491238396e-10 0 6.386467491238396e-10 0.00021 6.486467491238396e-10 0 6.486467491238397e-10 0 6.586467491238396e-10 0.00021 6.686467491238396e-10 0 6.686467491238397e-10 0 6.786467491238397e-10 0.00021 6.886467491238396e-10 0 6.886467491238397e-10 0 6.986467491238397e-10 0.00021 7.086467491238397e-10 0 )
X66 SYNAPSE 65 64 66
X68 CONFLU 57 0 0 0 68
X67 CONFLU 55 60 63 66 67
X69 NEURON 67 68 69
.temp 4.2
    .model jmitll jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.15mA)
    .tran 0.008 500p 0 0.008p
    .print PHASE 36 0
.print PHASE 52 0
.print PHASE 69 0
.print PHASE 23 0
.print PHASE 26 0
.print PHASE 28 0
.print PHASE 30 0
.print PHASE 33 0
.print PHASE 55 0
.print PHASE 57 0
.print PHASE 60 0
.print PHASE 63 0
.print PHASE 66 0
.print PHASE 39 0
.print PHASE 41 0
.print PHASE 44 0
.print PHASE 46 0
.print PHASE 49 0
.print PHASE 6 0
.print PHASE 7 0
.print PHASE 8 0
.print PHASE 9 0
.end